version https://git-lfs.github.com/spec/v1
oid sha256:1b7324883ed9236aa7a2987e45387e58f99d9508a83529e04b1c0569a7c50d00
size 13489
