version https://git-lfs.github.com/spec/v1
oid sha256:cb319f1d6abb8aa24ac697ee239996e0ef1731b7eb8f872b1cc1d687f64b4c36
size 855
