version https://git-lfs.github.com/spec/v1
oid sha256:918d6e5eea7de19322e15fc6b73d72fd6a3645712bae2afaac2e79909d30062e
size 845878812
