version https://git-lfs.github.com/spec/v1
oid sha256:3e41a409eaaa6cb33353022009021dccd6d7a6a7803632f76a1453d1790b3a39
size 67317985
