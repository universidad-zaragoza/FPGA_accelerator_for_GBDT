version https://git-lfs.github.com/spec/v1
oid sha256:e5b1bc014fb6b0ab317b0b4c6994dfc047cd4d1cdf36f68dfd011d7afc3ccc37
size 605
