version https://git-lfs.github.com/spec/v1
oid sha256:50065cdc37a40b54b9a6674397b1396d9d2197a7fe03123b11db0486945a5ae2
size 146439738
