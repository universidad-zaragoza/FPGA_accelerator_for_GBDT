version https://git-lfs.github.com/spec/v1
oid sha256:5326e47fe1ee0a18bb7463462d6044803d6e80ae7cfbd6b447188a9301a3cddf
size 764
