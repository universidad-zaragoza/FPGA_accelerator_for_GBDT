version https://git-lfs.github.com/spec/v1
oid sha256:8f13d71d93e235f791b38fc8a1264b010014f2a1eb6fdd1af3ee67eea1b1ee19
size 2335
