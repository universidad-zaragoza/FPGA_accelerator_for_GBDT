version https://git-lfs.github.com/spec/v1
oid sha256:105b90702257d421b2d10a56e8c8b7bc1625e171e907fff1e8d0730f86caaf1e
size 879
