version https://git-lfs.github.com/spec/v1
oid sha256:910f9138c3403828f65ed6381c3c17c237a713ada01e7e189278e46e2c1af38f
size 20571
