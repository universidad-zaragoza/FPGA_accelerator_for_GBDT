version https://git-lfs.github.com/spec/v1
oid sha256:43539c9e58d6d8d524cddb388a64923864babbaea50a7fa57e8e25abb5326e9f
size 935
