version https://git-lfs.github.com/spec/v1
oid sha256:73d7f24b969240e820cc519c8271ff9a8689f6d468be7ff1e4b145cc08c111cd
size 1330
