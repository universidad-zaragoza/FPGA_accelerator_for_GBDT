version https://git-lfs.github.com/spec/v1
oid sha256:53998d9b6042a448c02c2c608710509148a5605eac99fd2ed058e626b83b52dd
size 325482615
