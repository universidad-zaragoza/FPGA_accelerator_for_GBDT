version https://git-lfs.github.com/spec/v1
oid sha256:ad90860350e44301c69cffa4b584021fbfeb52ce5b8a5f57ab12cfc3c5761b10
size 16361
